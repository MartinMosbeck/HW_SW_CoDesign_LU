-- Load Altera libraries for this chip
library IEEE;
--LIBRARY MAXII;
use IEEE.STD_LOGIC_1164.all;
--USE MAXII.MAXII_COMPONENTS.ALL;
use ieee.numeric_std.all;
library work;
use work.audiocore_pkg.all;

entity audiocore_Simulation is
end audiocore_Simulation;

architecture testbench of audiocore_Simulation is
  
  signal clk: std_logic:='0';
  signal res: std_logic;
  
  signal Istart, Iend, Ivalid, Iready, Ostart, Oend, Ovalid, Oready: std_logic;
  signal Idata, Odata: std_logic_vector(31 downto 0);
  
  signal lready, rready, lvalid, rvalid : std_logic;
  signal ldata, rdata: std_logic_vector(31 downto 0);
  
  signal counter: integer:=30000;
  
  begin
    dut : entity work.audiocore
		port map
		(
		clk   => clk,
		res_n => res,
		
		-- stream input
		asin_data => Idata,
		asin_startofpacket => Istart,
		asin_endofpacket => Iend,
		asin_valid => Ivalid,
		asin_ready => Iready,

		-- stream output
		asout_data => Odata,
		asout_startofpacket => Ostart,
		asout_endofpacket => Oend,
		asout_valid => Ovalid,
		asout_ready => Oready,
		
		audiooutleft_data => ldata,
		audiooutleft_ready => lready,
		audiooutleft_valid => lvalid,
		
		audiooutright_data => rdata,
		audiooutright_ready => rready,
		audiooutright_valid => rvalid
	);
    
    stimulus : process is
      begin
		res <= '0'; wait for 20 ns;
		res <= '1'; wait for 20 ns;
		Ivalid <= '1';
		Oready <= '1';

		rready <= '1';
		lready <= '1';
		
		
Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"61bdc2a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1423a44";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57afd3c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc544d37";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b9baad3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d476651e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b828ae6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d7969118";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c4f6ad7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0afae37";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4d3149ae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1c4a952";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"583f57ad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6bdbb57";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5434529c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"babfbc68";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"59322f89";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a9ccd175";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6d25396e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"80d3e1a2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8e17264f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6cbfb7a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a5363b3e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"51beb6b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a44a5b44";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ea7b8aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ac472d53";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"60b3c2a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2513336";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"37acc3cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf5d472b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d96acd4";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"db5f5327";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"20849fdb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d48a651d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"0f7f91ca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ce837a3d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"27747ac8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d778733b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d9086bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"de7b9035";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1e6c67c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d87f9d3c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1c5246c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d8b7b33a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31523bb2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bbbacf57";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"453b23a6";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"9bb7ce79";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"683d1f7a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92cac37d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65443f87";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8bb5d079";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72421f93";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81cacd73";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d36206f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5acae19d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a3372f68";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"37c6cdba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d6453b4b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"33b4a5bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d1695540";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1c9795c2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b76f6b53";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3e9e8bbe";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d564733d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"34a68bc6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d36d8b36";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1b7f66d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d28f9a31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"27693ed3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dab9d447";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"304e2cb0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"abc7e475";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"613c209a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9cbcc782";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82453875";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7fc8de88";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8c46337f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"69c2d39f";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"a93f2165";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4fc4ceb2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd5a3845";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2faecad4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d05f633d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e8f98c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"f67d6e2c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"207184cf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0979b3c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31766dc9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf9b924d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4d7168b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d087993b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"27776db8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d199a741";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c6250d2";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"d79eb936";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c553fbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cab2e83c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"49462fa9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5bfdb6b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"682f3195";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9cbfc363";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7249448f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85bec85d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6f3732a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8fbdd05e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a292789";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74d7e275";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9a30316e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50d5d59c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc1d3450";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"2fb3b3b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dc4f5e27";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"169f95c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc6a7b45";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"368572c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3718239";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"32857eb2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd7a8939";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"29786fcb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd748f2b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f6a49cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cea1c125";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"374e36b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bcb5e047";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5a272a9d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a5bbc15e";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"73443495";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7dc5cf5a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f39358c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7cb4d472";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a342684";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6eccd079";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9d313e65";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4bd5cca0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d233474a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38b2bcc2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"f6586e29";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"198786c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc7c8e32";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"226556c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d6959f45";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"405750a4";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"bcb8c255";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b464594";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9dacbd70";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"66362a8d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97b4ce74";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76442672";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"80c8e688";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"89342357";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5cb5c9b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b53a2a37";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3dafbbba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc604f31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31949bce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf735a4d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"46868eb6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b27c6240";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"459d97a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba525a4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1f909ec1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d1586136";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1f998ecd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e27e8131";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1b7466d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"df87a73d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"295854b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"caaea33e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"395f50aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aea4b65f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"484842b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adacbd59";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5d5a36a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1c4dd52";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"60392da1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92c3e782";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83290a6f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"59d2d29d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b64d3750";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"36acc9c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb614f48";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d97a6c2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc70603d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4192a2b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd717240";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"308293c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e8707341";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"287f8ac2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd95992d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"22675dcf";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"ea8eb639";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b4d49b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dbb5d53e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"46423e9b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aabdc86d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6032399a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9dbbc274";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"793e327c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"90c1e06f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"803e3e73";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7abbd496";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"91331e60";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5cc2d098";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7452a35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31a9c1d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d36d5732";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"1b708de4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d9978833";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"30625cba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bdc7b043";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"444055ad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a3b9af72";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6a414e99";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2ccb26c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71494588";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96c6ca7a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"69324b7f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"98c6cd90";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82292b5b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81d7d2a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9e2e3d46";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ecccdcc";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b0444835";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"55a6acc5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b85c5336";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"56a1b0a8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6565954";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"499dbaba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2504240";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ca1c2c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d16b4a2c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a8ca2cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"da766a2f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"157172d0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d39b803f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b626cc0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6b29d49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"384865b7";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c499a144";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c533eb1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfbdb351";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"354936a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3d5c670";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4f2e298c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"99d8d083";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75222763";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74d5d9aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85381e4a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"52bfc7ca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af533c3a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48b0afce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b15d593c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"439d9dc2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b25d4f4a";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"49939fc7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c081652f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b8ea2c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d477692a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1e666ddc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d9a2903a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"244c50cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cee2b94b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"442c41a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94d9c678";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77213978";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8cc8bf89";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"793b4769";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72d0c5a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8b3a3f66";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"73cbbaa5";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"ac364547";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5abbc5bb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7564f35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"339da5d8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c96d7021";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e7d6ee3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d191a81a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"395959bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"afb0c653";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5c403fac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9ac4a769";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7959458f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86b0bb56";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"603b48a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86cbba76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7d252d93";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"7bebc384";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a2e476e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5edec19d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1214a52";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54cba6b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8475c47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4fc2aabb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6526349";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4daca3bb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ab4a5449";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"53aa97c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2655829";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"35ad9fd9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4637a29";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42897eeb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d185981d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3c6d67c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfb3b332";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"474845d3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aec0bd47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6d3943aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9cc9c048";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"673b4c8e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82baba71";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7a2c439d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"95dbbd6c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85234276";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fe0d28a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"930c354d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57c7aeb1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be224b2e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2ac19ad3";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c15b7529";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"279d77d7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"db708c30";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a7a6bbf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0899532";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b766bbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b28a913c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d6452d0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c29aa534";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"49513cb5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97c5d43d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"612821b0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71dbc779";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9a2f1680";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"47d9d49b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf454952";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"30a9acc3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca5e5249";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40a695bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7706d4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31988eb8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c37e814d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b7c71cc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e18f9f33";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a6857bb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6acc752";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"344834a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bbc9d869";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"723f3386";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96d1de7d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"87322b5c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"63afdea2";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"9848315c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68b3b7a1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a0514d5d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"62b0c793";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a4464b60";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"52a5c6a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1463153";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ab5bcb9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c65c4e35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1f92acd0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d76a6a31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e827ec1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e28c8436";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a787ebb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc898947";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"357467c5";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c57e8743";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b7e62b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c684ad39";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1f6d4bc0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5aebd4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"434624bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b6cae064";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"593f159d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86cef386";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92362772";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72c7c6a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"99464059";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61becc9a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2464871";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"60b4bf9e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2463060";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"53bec4a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be434658";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"32b2b9be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd585534";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1b9787cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ff7e9125";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"275d78c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d299953f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38615cb6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc92a949";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"386652b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfa3c344";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c4a46a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bcb7d65b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5c372593";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"99cdeb70";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"6e362075";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ebfec96";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b2c1e51";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"62bbd9b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ae424836";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"43adbbbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd59673e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"418a9bc0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd765c38";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42888fbd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf807647";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c7d8bc3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d8808632";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f6968b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d7959732";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1b4253be";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c7bec24d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"303234a1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9cdc765";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"64302981";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8fc9bc72";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58384494";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"95b9bf70";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"654d2d9c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9dbcd15f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54461f94";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86bcda70";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6d340b8b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72d8e08f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a32e106d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54c1db95";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a83c2e5b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"48bcc1ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3543d6a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"59bdbf9f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af464567";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44bfbba2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb3c4359";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38c4a9b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca4e473d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"21c19fd2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e6617b31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"168f79d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3728538";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b8664cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8909442";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b7e71c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8859631";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"39724bce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be8e9b20";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"326743cc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"afa6ad3c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"434734d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1c2c345";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5e3431a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82ced855";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7a2b2387";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"78d2c384";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8c3f258e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"60cbbc86";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b473e78";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57ccba89";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"93343776";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4bc4b1a4";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"bb3a434e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41d2c2b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf495a3c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"27b08fd0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d35b7d2d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1d8c64dc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d785932f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e8058c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c79aa845";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"456557c2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b58fa543";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"416a59c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4a6ae34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"46604bd9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0add146";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"593534be";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"a4cbd54d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"79341a99";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75e1e878";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"98263087";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65cdd18d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ab304d7d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"73d0b788";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9944417c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61ccc090";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8c2c3c6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75dbc997";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ab263b56";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"63e1c7b0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5214e47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ec7b4d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6435031";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"4bbca0bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc4c652a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54a3b3c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aa55603f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44aaa8ce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb595a24";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e9eabe8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc707216";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"327693e9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d08f871b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44746de2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cca79d31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c5a64c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"beb3a03d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e415cbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9bb964f";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"4e5461b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bbbbbe50";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a4759bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6c2b74e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e302c9d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bdddcc6f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5a1f398b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"87ebd696";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7b2a2f69";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83d8d197";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96393f52";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6dbebeb2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"904d4775";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6bbebfa5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a44a295f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5dc3c8bb";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"ac43303f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"33b1bfd4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1674434";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"32979ce4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e48a7526";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"257279da";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"caa59b35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"33485fc8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1c4924b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b5765b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b6c1aa5a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"435957b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3bcb356";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c3c2fa2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2dbc568";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5532358b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"96ede78d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76232b76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ececaaa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"982a2d46";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61d3c9c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"964d5056";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"63bcc2ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a346325f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"66c4cfab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aa4a365c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3fc1debb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba4a3d4b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45aabcd4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d75f4839";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2da6b0c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d36a663f";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"28999bc9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e1766243";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b8895bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf797243";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"249b8ec5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0717a4e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"29957ecd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e2748d32";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"218969c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d39cac3a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a613dd0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dcabc44a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"464b40b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8b9d74e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c5045ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1a7b359";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"68533dbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aebbc949";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"565132b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92c8da61";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6a3118ae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86d2d576";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d311e85";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"59e5e38e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ab2c2e68";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40c9b7a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5433e60";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3eb9af9e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aa51585d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40b8b2a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc3d4b4c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3fae97b8";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"bd4b5638";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"18b292cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d55a772e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b9369dc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"df839e1a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"255944d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"baa6bc48";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e593dc0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aba9bd54";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5c533faa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"afaebb48";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"524735b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92d4c25e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"66362aa3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ccfd47a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85351c78";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"65d3d08e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"99332960";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44d2cbaf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3413e5f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"47c3ada4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5495056";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"34afa1b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a456584d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42ae9bbf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c24c5b45";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3cba9cb9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc566423";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"27af94e4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d15f6d29";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a9280ed";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d78b9c21";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"31825edb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd90973f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d6c67dc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c198882b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"477778c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb958227";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f6f72e8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd999433";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"345452dd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3ccb327";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"423f51c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bbd2c651";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"53243daf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a3d3bb5d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6937478c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94d0ba70";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"602e4c92";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a8c1c078";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6c293487";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1dfce6f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"70263576";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"80d2dfa3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a132552";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6ecfcaab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a534392c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45c8bed0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b347503b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a9c99be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3695341";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b9aaab8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ae6b5233";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e92b5d7";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"d3665421";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a727fcd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c79a760c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1f5a6ccf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0ac9a45";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f4057bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5bda746";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4d3c48a8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"abcbae60";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a37539d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2b7c773";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5037408c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a4cfb973";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"692f2f7a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8fd2d68b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6b2b2672";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"79ccd8b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94312140";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ad0b5ba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9e493e42";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3db9becd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba504b4d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45a3a0c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be6e4e41";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ca6b5be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ab5d4b41";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ba8b1c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d5563c36";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1a93a1dc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"df8e712e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"0a7a8fdb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e3a99536";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"2f5e61c2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dda99e4c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"305e5bb7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cba9af52";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31706bbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d2929740";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"376955c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dc96bd3b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"315a3fc8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"deb7e538";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"444c35b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bcb6ce5b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5c3a25a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9abdd256";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6d4a3e99";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"95b2bf5b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"683e47aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aab1c14e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5d4c38a2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9cdada50";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"771e3090";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76cfe57a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97193178";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68cec67e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1423763";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57c4c79b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ab264b61";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5eb8ad9d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6354a4d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57d3b5a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b43d5347";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41a8b4d0";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c3365226";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38ad8cce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c75f751d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"338274dc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c97e9c20";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d6d59d3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb959337";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"476259c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2aeb141";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b564eb4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0a5b63e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"544d3ec7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0bbb343";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c2f3bc3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9fe7d04c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"601633a9";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"8adfc974";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"981b1c87";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71f7ce90";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9432516e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65ccbc98";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9434486d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82c9b699";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"923b436f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ed8d99a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8b333d5b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6acec9b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b62b3038";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"53cbc0d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be445d25";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"43aab8c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be615929";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"478d95c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5645f3d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b95b2b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb685e2f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4293b8bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d6614934";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1991a2cf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e074641e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1b6a89ce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d99b8424";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"265d70be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc788f41";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d6d77b0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0987c47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"287585bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d2778837";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"1a746ac7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e07c992c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b7649ce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d093ba42";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1b5d3ab9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5a1be44";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"404c2fb0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aeb3b744";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"574e4cb4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9faab956";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54553fb3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7aaad3e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"533f3bb0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97c0bb4e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5b3239aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85d4d15e";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"872d148b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"69cfc67c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"902a336d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3bc8c29e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b4c476b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6ab7a392";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9d444a6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5dc7b497";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8936415a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5fc6bcb0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a72e353c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5bc3a7d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c545621d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"16b190e2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca658129";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"288d5cda";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"d3899329";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"437767d0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af95993f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"477378d7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9907f36";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"457262d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5aaa030";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"28546bd4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9c0b039";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"442938d6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2dbc047";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"67283fa4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cfa09f34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"394062c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cbb59a51";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4f4c5b9f";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b2b7ae51";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"484f4ab2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4aab359";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"434239a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bdc9d160";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4f362882";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94d2ce79";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"671e1d89";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"79d8d9a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8537286d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fd4d39d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b473158";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"64bcbfa7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d42316f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"59bec99e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a8483265";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"5dc1c5a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b546315b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2eb5cacc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c655444f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2cb6acc8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"db654c38";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1fa59bc8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca736e40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"268885c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d77b7142";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e9b86be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd718d39";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"208d71d0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dc7da23f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b6c47cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dba9b942";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3a5444ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"afbfd45d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"573d20a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9fc6de6c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86452781";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7cc5dc8d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"873e3974";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6cbcd799";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0472a6c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4cbec6ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf515352";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"903f3760";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"53bbcc93";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a53b2d63";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41b8bcab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba4c3e4c";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"44b0bca2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c752543f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"34969eba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e6546f38";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"0c8476c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e08c942e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"215f56bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cdaeb946";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c323c9e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adb7c75c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6b412686";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"89cac17d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6f444172";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76babea0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a393866";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72b7c190";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"9a453549";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"55b8ccaa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ab484638";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d98addc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d46a5f16";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f8491c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc8a8030";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"324e72cc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfa79f3c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b4459b0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3bcab4c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"56464cae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"98c5b466";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57364e95";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9bceb078";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6831337d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"94d0c27a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f273b67";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61d1d0ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"90313b46";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"52bbabc6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf474e2f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48b097c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1616d41";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3aa1a0cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc62523d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54978cc8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9767026";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"308381df";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8888239";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"33716ad7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d5a4812b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"35535fbe";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7bea437";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"393954b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adc2ac63";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5d4037a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9ad0c46b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6b3c487d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7fcdb98d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6e363879";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7dcdb08f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8c38486c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"67d5c6a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"90373e42";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50c8a3d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be3e4625";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"35af88e9";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c76f8a2c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"288b68d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9909137";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"466454d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3a3953d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c5a59b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a69fa441";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a4d53b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7ab9857";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"59413baa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"90d9cd54";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6f203789";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"64cbc884";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7242a63";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40cdb0af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1584e46";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"30b695c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc647545";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1b8a6bbe";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7808d49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"386b55b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b796a845";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4063509f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9ea6b654";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"514b30a1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adb4be70";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"653d3077";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77c1da8b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8b37305a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"52abbdaa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4563549";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"409aaac7";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"bf7d5f35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"357e92be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b77c813e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"426b7cc1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd90813f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45656eaf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5949137";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"334f5fb8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3a0a44a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"434855af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cbb5c146";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3247409b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4babc65";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5a2f2ea0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7b8ce71";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"73353961";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"83c2d385";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82494972";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76bcb992";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8f323a6c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7eb4c98f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9e4a3d49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5cb8cdb3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b54f4738";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b89a9d9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d275691e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b817fcc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb91912b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"32485fce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3b8a943";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"583b549c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2c9b44f";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"5a3c4a9b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8eb4b370";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"70294290";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9ecac677";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"732e466b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7dccbe88";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8e263f5d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65ceb9b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6264739";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"55bbc1be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba546323";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b9f8ed4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf627f2f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b7672c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf929432";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d7178ba";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"ad96933e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50535aca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aeaeb636";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6e3f3fa3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"90bfcd63";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81313387";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6bc1c589";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a8324369";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ebdb9a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c84f6040";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c9f9bb5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf677748";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"37836cbb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d575993e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"386c5d9e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2a1b654";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"535350a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1a8b263";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5e52499d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adadd75b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6547348b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"93b6e173";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"773f2b81";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"84c8d68e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"953a2465";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"60bad395";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a647425a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"55a9c5aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b04a4d6a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fb5b68a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a0514d6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57b5c09b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b23a506d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4fbdb7ae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d746523b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31b9a6b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd5d763e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"28897ad1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e67d983f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a7167b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb9eac4d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b5c4db0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cba0c05c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5e543ea9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adb4c960";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"604c3795";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96bbe181";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7a46278f";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"83cce795";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b3d2465";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58cbd2b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a84c4050";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"46b0b7d3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4634f4c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42a1a6af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c56e553c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"29a09fbe";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc6c6750";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c888dc8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e27b753c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1f9e7dc4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3949640";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"26684fcf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dba3af43";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"2c544cad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3bdbc56";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"424c37ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a8c0cc7b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"643e2283";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8bc4c68f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"753d3d5e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6cc1bd99";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8e493d6c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61acbeae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ae58274b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3caeb1c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a66c5234";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"338193ea";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"db8d752d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e6267cb";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b9b6a531";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"393755bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"acd1b252";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"762d3ea2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"98ceb56d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"683f468b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8bd2bb76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6b404795";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a4c8ba77";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6c2c3b81";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97dfd481";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6b373573";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83d9e09a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f222d76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"89c8cfa0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8b3a3756";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"6ecfd090";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a413477";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fbacd9f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"933e1d6b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"69cfdd93";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9a46305e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ac2dbb3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb3c375c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31b3b3c2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd6e4c2c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1d9ca7c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"da7b754b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"36797bc8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"da8f8d3b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"288169bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"caa79f48";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"335459c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d1a9b74c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"434d46af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bec6c758";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"414629a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"accfd780";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"563d238e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97c5cf81";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"743d2576";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77cdcd95";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86441c83";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74becc91";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"814c2579";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76bcbb82";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83412b7e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"64d0d08c";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"9c36246e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"49c9d0a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd422a3d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"21bcbebc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ce52573b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"248e98cc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e06d6e39";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1d877eb9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf7f843c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c7372c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5849447";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c705ebf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cca0bb35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e5e35b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bca9c75a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d341c9c";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"a3c7d470";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77352073";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ec8ef86";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"87341663";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"63c1cab5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9a4e2856";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58b9c1a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a852435a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"53b1c09b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6412861";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48bdbf9f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b549354e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"36bcc0aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf3f3e42";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1fb0a4bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c64c5644";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"35aea8b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7526142";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"35a49db7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd41583c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3cb89ac1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf536933";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2dac98cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ce607a2d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a8776d9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4778421";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"307b57d7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c282a72b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a6e59c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3a1b83f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c5d44c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a8ab9e3b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"4e565dc4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7b5ad47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"51504ebd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1bbb73a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"533136b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9ae3c465";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"602936a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7bebca76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"921f2d78";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72d4bd89";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"913c456e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ac6b4a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d414166";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"73c5ba9a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94333e5c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ec8c5aa";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"93314044";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ac2abd1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc4f4426";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44a999d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c35e6f26";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"328b81d8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba75732a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b7e71d6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c199822e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b6383c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b69a8e32";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"354e56c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7a69332";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b4448b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0cbc245";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"462148a5";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"a5d4ba60";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6a0f2588";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7de9c57a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82233c6f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5dd0c19e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"931a3c5d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77ceb995";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"992f4248";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"62d4c8af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97294746";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54b7c1bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc373f27";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48bca9c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b44b4c24";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ca3a0de";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be55572e";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"439b99c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb6f6825";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3683a6cc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be736f3e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"418397c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca74602a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"328790bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d2797c2d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"126786d3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e49b7f33";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a6360bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cbaaa63b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"234e5bbf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2a2ae49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a5752ad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7a3ab51";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"405b57a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c69eb743";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"374d3db5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6adc946";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"584e29a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aacbee6c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5e2e238c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8eb8e07a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7e33167d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81c8d783";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96443b78";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6cb8dc92";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6433774";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6dc0c78d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ae48385e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4dc9d5ae";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c7394f5d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"34b9b5b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"db59493b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"26aa9dc5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"db6a783e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1d8b7fde";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d791893d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"35886abd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d48c9d42";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a7263c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c884a33c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d5f40c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4b3b13e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"49563fb7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9fb6cb5b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a3d1aac";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"9dbdd35c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74371d83";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76d1d185";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7d323289";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71bbc77b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9a413169";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61c5be80";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97403674";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"59b5c49d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2394163";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54c9c298";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c536324b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1ebab5b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd33543f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"24ad9aca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dc60662d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"2ba383c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d4637f3e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b9081c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c65e7c2d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"399587c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7658129";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45948ed8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf668612";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e7f62db";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca8ca412";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f5c53db";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3a2b12b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"52445dbd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bbaaab2c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"515659c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1afad47";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"47475ec4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6b3ac3c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"534c54b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bcc7bc43";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a2148b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"add1c167";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7425328f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92e8d27b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6e3e4285";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8ad1c399";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8b25456c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"80d2be92";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8350436a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fd0c2a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97363463";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"62cabec5";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"a93f4d31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42c2b0c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b35b4f38";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c9d99e8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c66d623f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"32919ac5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c27c7423";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"39767ad9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c486783d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d7371d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfa89837";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d7066c2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3a59e41";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"323c45b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"babfb74a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"372933a9";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"9aeecc75";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"67302987";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88dfbc9b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8b223663";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"69e1c2a1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86404a62";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5cc3abac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1453665";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6db6c5ad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"984b3f41";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48c5bcca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5553c34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44afa6ea";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca6a6333";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f95a0db";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c87f7022";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"397883de";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d1967237";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"39727cd6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b699913c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"317476c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d7948943";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e6572cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cbaba13f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"294657c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d2c9b749";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a4036ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0cdc469";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4433388c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9dcdd477";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"603c2c8e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96c8c083";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"74363f87";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8dbfd570";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61451698";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85d0cf88";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8639106f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6cd0dba6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"933d345f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50c1c5a1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2462954";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48b5bab4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b556444a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"339ab5bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2614f44";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"379891bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d5746033";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"13868dc4";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c9777c3e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1c6a6ec1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e3929430";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"21584eb4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c9a5c343";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e3033aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bcbccc5f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"59322574";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96d5d487";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6a283974";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72b6c089";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"89432b6c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7dc1c58e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8b434357";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68bad9b1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aa35333c";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"4eabbeb4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca5b4721";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b92a6dc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d27b752b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c5877d9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0ad921e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42506ab6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4b2ae4d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c4b5db3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bdada75c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"53454ea6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9c3bf4c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"554148a6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adb7cb6a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5d2d318c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3d3df80";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"762e3068";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7fe0d4a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"95283c65";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6bc4c5ae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2434543";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54babfac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a5534157";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5aa9bdc0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5514e47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4dafbfbf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c25f5335";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3699aad2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dc726432";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d8198db";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d68f8128";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f7388c7";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"dc8e893d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"33656bc4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dca19540";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"24616ac5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0ab8f4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b6b5fc8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d2a1a644";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"296152b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6c5cc5b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"37432aa9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6d4d678";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"66332f83";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"91deee8c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7c302d72";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"73c5c9a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"99422856";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"67c0cb9a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d504263";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5eb3c8a1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b142385f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4eb9beaf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c24d373e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"24aca8cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb5f4134";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1a9093d7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d98b7832";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1e7d75cf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd939739";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"275760bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6a79048";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a5d5fac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7a2a156";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3d4c49af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d5b3cb4c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4545388f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a4c6d871";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4f221588";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"89c9ce8c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"872c1e5e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65d5dba5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9e473e4e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4faabec3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b747393f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50a0aa9e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ae5a4c46";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40a3c5cf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2574d46";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c99aec3";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"da6e5921";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d8ca3bb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"db5f752d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"227d86c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e0788234";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d8282bb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd8a8c3b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"316577c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d17a8734";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e8070bb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3809835";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"277f68d7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"df83a735";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"356552c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3a5be1e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e5747c8";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"bca6c940";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e4b2bb4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"acb1c24b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5f5355ad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a3b7bd42";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"60414abf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0aeb045";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"544a47bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1cfd450";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"643738ae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9de0cd68";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81183588";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ed9cc7e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a23437b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fcaba96";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a84c4472";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"7ccdc395";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7e414373";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77d2c39c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"912e2d5c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6ed6c1ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9737444b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4acbd5c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1414349";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ab7a1cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b253512c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42a9aabd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a15d5446";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e97a6b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b75d4a40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"419baab3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5634f34";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"2794a5d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d6726830";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e737ccd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d89b892f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"245567bb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c99d9139";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d455eb1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bdb0ab4d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"384e53b1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3b0c153";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4d3f409e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1bbbd59";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"43343397";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"abc5d46f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"62352d91";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aed9ed70";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"77322878";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8ac8ed83";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77373782";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85bfc790";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"874e3989";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"87c2ce6a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"754746a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8dbfca6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72342aa0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8be5c76e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81312a8b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fe0d881";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a28388b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6dd3bf7c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94443979";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"66c7bb82";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"76354c87";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"87c4b077";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"78253783";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8fcfc977";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"761e3b72";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75dcc6a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83362461";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ecbc5a6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8c394150";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65b9c1a6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8f3b3663";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72b3bc8a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"91483d64";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"66b8d393";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9c463067";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5aaecea7";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b840333c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48b2c0a8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c04c4c46";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c91acb3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c55c5a40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"509bb0ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc615f51";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4794abb1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba48594f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3cb8a0af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d45a6848";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3aab9fc7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d451703f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d928fb6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc6f6f34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ca588c4";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b96b8545";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f927dd0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1707937";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"46927dc9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4848f31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d7b72e7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc869b35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"476851e3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1cabd31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b4944c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a8c8cf57";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"712641b1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"89cec165";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7d403e8f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83cdb878";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f3b4a9d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"98c5c26a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74394484";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8de0bf76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68283296";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82e4c78a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7b312d7a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7aeace8b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8731476c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72bfbb9c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"782e3470";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88c9b17c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"744e347c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"80c1d777";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6e36258b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8cbad976";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7a341676";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"77c5d779";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85372a7d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"69c4c18a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8e3c397c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71c1c677";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a414580";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77afb77a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88354188";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82ddc57c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9a3b3f70";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5fdad19e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b925496b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5abfb4a1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b84f5648";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"53c5b4b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a4515b5d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"65aeb1c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b747593f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58bf9fbf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b64f6545";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"43a8a6c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b85e5838";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44a6a0c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3706432";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"398b94da";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4716826";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"408483bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3806c48";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"478ca4c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c26b5b52";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a869cb7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ce735534";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"2894a6c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd777e3f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c7f80da";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ed989138";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31686ebc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bcbca852";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b5355b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1a7a660";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e624ea9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9bcbc54";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5455499e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a3b1c06c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"513420a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9dcdd470";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6c361f77";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74d3e399";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"912f1d5a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"63b8cba8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a54b284e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54b8cfa6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a14a4459";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"62b5be9e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a33b3a61";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58bdc27d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a53a2e66";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"47c1ca99";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b020395e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50ccc79e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb2c454f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"51c1b79d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af344b6b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"64c3b195";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"9938435d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76cbca9a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"91284266";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7fc7c2a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a0304b49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68d0c3b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96444850";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58b3bebd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a740454f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"69b1baaf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9f5f5248";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58aabab6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b34e415a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5aa9b8b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd645c47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2eada3c1";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c9644d37";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"307e87d0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d37a6e2c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"166e7bc9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c884843d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"375c68b0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf918948";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"397377a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c57a8b40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"347577c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d97d9336";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38816cd2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d694b53c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"34755fc7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d090af3e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41653fbc";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"bdb3b351";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b635ec8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ac9aa247";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54684fb9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2a6ab34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3f4c4dcb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2b5bd50";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5b4235ba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a0d7c05a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76362e9c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6bd2d97d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9a242d80";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"52caba9d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2463258";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ad1bca6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a849535d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"4aafa8b1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb475045";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4bb9a0b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd4a5a3e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"23be94dd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb62693d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"37a078d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb67821b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"308f79ce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be6a792e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"378b83d8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3776e2e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e8993dd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c074701c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f7c7bda";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c8786a2c";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"307b83d5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca957726";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"296983d6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d8968225";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"345970bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfa48d36";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e6273be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba82884c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"376870b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e5a19738";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"246261b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0a4af40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e4b42b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"beaebc40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a4c2ca4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adbbd066";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"52322c9a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8eb5d36f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75432b70";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"91b6c46a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"72363183";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86bcd275";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"843d3979";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"78c3dc77";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"93312e71";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65b9d9a6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b83b2a58";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"43c4c9ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c14e4d4c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"36aeb7ba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d94e5a4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4fa39fad";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c86a6644";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2da2a2bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc647057";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"36a586c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd6f8636";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a967ecc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf90a036";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"236845d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d5a7b545";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"465a36b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3bad758";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b4434a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9fb4cf6b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"70411e8f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8ac3cb70";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"723d2984";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"60ccd084";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9933226a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ac2c298";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b446294d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2db8bcb2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c74b4d49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2fa6a6c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e2625832";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1b8f8ebb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d4787e43";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c7585bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d476803f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a8571b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d2799936";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f787fbe";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d37b9d35";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"2c7357d0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"eaa2b03d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"376150d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"beb6de4d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"484731b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5bcca54";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"634c2da3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"99c1cf6e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"674943ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97bbbe62";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7444329b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8cc6c85e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6c28289f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75d7d975";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"982e2271";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"56e6c884";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"992a3a6a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"43c8b1ae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc314352";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3fc2abaf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc5d594e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3aab9fbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b6476148";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"39a687be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c15b701c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"26a77cd3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf6b8e31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"29795ddd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d58eac1d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"325f47b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9a1c23b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4f422fb6";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"a3aec856";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6a452c8c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"91c3dd5c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76373f9a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85bec873";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"98252986";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"60d0d27f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af3f3a5b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42bac8a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ce354a51";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d9ca3af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d9506d2f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1a9a98c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e7738f32";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"30685fc8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e598a740";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3d5b5eab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4b0b452";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41584cad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bea2b154";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"514d3cb1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"acbec65a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50452b9a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94cccd7e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7b3e1889";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7dd0e095";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"91462567";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4dbcd3a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ac48374e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4baaa8b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9564856";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41a6b6aa";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"af635552";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c9ba4b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2585246";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"369e9bc3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d36f783a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"17918bc9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e87b8337";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"206d59be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dc989f37";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"24625ac2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfa1b654";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e4d3fa6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c49ab24b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"405746a6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0a0c74a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b5045bf";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b4aec843";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6a402ba4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9fc5ef57";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6e322883";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7cbecf74";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92372376";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"70cdd68e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1385078";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ebdd0a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b24a3a60";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5dc1b59e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c9524549";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2ebdbdc3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d254654a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2aa49ac5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"f07c713d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"259287ce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d7789b34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"206b62d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e4aab341";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a613db0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9b9cc58";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44543fae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"abaabc67";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5a493097";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2c8c861";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65443497";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"87bacf72";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77320989";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6ed4ce7a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8f382150";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ac2d7bb";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"bd3d3951";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"379ca1b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca6a562b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1b929abc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c57c714c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b7282c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0837b3e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"217b73b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca878841";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1d7564c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dc8ba142";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b5451b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d1abc940";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e4d2db1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3aec65a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c412a9a";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b0b8c65f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5d453791";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92bcd760";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"703f319b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92b8cd63";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"723f2d91";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94beda52";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"772b3187";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"70cad983";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a52b2e78";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"64cacd81";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9f333160";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57b9cb98";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a23d426b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"63c4bc9d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7364f54";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"53c1b7a8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a82b4259";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ec0b7b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb3e5438";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4eceaacc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0456d25";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2fac8dda";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb647935";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"35a280db";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c8818631";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d8075d9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b17b8132";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"467f77d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c687822a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a7d70d9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd8f9a25";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"385658d5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8ac9822";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"414145c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1c6c63c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"582642a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a3c2c359";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"78324495";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"93c9bc61";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6f38589b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a0cbbb79";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6f313890";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9addc286";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"70363f74";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85e1d99f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"921d3457";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6bd1b8ba";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"ab284439";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ad5add6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af595445";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"43a68fd8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b85c5c2b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"489b9aca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b06d622d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"399395dc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c9695e26";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"328692d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ce8a6f10";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"196277ef";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c69e8627";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e4d5ed7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3a59237";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"346976b9";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c2ab9a30";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b4d5cc3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d49a9c45";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b595ab6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ccb2bd39";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b4949b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7a2c04e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"403831a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cabdc64a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"534b49a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"acc6e067";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"603e2e9c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aab6c164";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6355439e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a5b3d357";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"574c41b6";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"abc2c94e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"663922b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8ecadf5f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6c3f289c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"84d6d473";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"89333194";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83c8be6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75324e8a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7cd0b67a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"723b3aa1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8ec8b97a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6c413d89";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81d9c97e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6e202c74";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77d1b79d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b1c3c56";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"5bcec0a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b3f4a4a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61b3a8b1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a63f534b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"60a7a9ad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a3565143";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57b6beb8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aa4d494b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"509fbfc9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc5c501b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"388da7c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c47a7929";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e758bdf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d090893b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"406d7ec6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8a28d3f";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"355e80ba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4998043";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"365170c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d8a5a03d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b5e60be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cabbbd4d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"414740ba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ccc4b260";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"454b40aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bbd3c764";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e4a43a2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"abb2c967";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58392da4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7bdc659";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"485733a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a5c0ca63";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"60431dbd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97bed25c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"66340991";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6ed5d76f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"80372178";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6ac1d791";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a335347b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ec1c27f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96453a72";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5abeb48b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97353b86";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"67d0c67f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92253664";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"53dfbda9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af1b3a56";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4cd3adaf";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"ac3f4b4e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ac4afa6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ac455152";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"55acaca8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"903e4354";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6dc3c09d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9340454d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68b8c9ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97322553";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ab7c4ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a645373f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58b3cab8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b54e4d4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"559db3ae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b65d3953";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4cb6b8a1";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"ad5d5d56";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45a1c7b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c84a4b52";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40aba7b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d56b6134";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1a9390cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e4798941";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38656bc3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d49c9e36";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"326c6bb3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4a1a64e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"335f52c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6a0b143";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"476144a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"acb2c154";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c492fae";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"afb9d372";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"643f1c9c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"93cad960";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"733c278b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75c9d081";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"87351b87";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71bac287";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8e4e3a76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"67bfc579";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8b3a3d81";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"70c0bd84";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"95283182";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68dcd07e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a22f3365";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50ccc1a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2203b53";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"49cfafac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba40563c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3cc5a3b1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2496356";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48a39fb9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a24a563c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4fbda7c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b74e5929";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38a597dc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c9496f18";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b8679d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ce828e0a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"307f73d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3888e34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"435c69d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be9a8f31";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"38706cb4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba988c38";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c5a7ad0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf8b8a27";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"365e72c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"daba9932";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"274c66ca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cea6ad47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"394d58b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0b5a447";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e5c61a2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c19fad54";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"385753b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cfa4af4c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4d6642be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5b5c84b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3a593bb6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aeb7c55f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"613d2aa0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9cbecc64";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68473794";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8cc3df7c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7645218f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"78bccc84";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"914c2e6b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61bcc784";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d403178";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57c5c6a6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba44395f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3bc4b3ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca4e4f43";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1ea69bca";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"d2686d3f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"228f7ecd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d98f8d40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"26836ac7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c9859043";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"376e60b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3949a49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"387561c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c09aa947";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"336545c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c39ebc37";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"384825af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a8bcc952";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4d3e24a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97cacf6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"713f1b9d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"7dc4d062";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"813c278c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71c2cc78";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"823a2a8d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7bc6cd7b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8f352a78";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ed3c789";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94262c6c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45d3bfa8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9404153";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"34c1b0b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cf4c5d47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2fbb9bc4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc536745";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40a591bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7636747";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"31b692d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb597b3a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a9783da";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c272731d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"33907dd1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd7e912e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"377570de";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4929132";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"446d6ad3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5a68b27";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38627fdf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1a29836";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"405b68d9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c8b69d38";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"425563c2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7bcb443";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3d3748bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"baddbd57";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"642937a1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9cf2cd73";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71293f88";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81d6c094";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f2c3d76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"80d2c194";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81434b5d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"78cfc6aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d2a3e5d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6acdc3bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7463d36";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"51c3bed6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba515f2d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"388fa8e7";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"d66c7a1c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c8b6ee1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd949f2e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c6674df";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0a79043";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e5b66c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3b99d2d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"47505cc5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"afb3b354";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c2e3fb6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7d7c259";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"612c418d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9bf3c776";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"731d308a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75e0cba2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"942f3f5d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"58d6beae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b34c5342";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ebbb3bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"993a504c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"52bcb1c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2544b35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40b5a7cf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0585f2e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38919ee5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd756d2e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d8f84dd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c98a8526";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42747eda";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2969137";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"305c6ed3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4ab8a35";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"406a65c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cba59d40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f5a69c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c8aaa03c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"354847b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cad1b34f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"393c47b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7dec768";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"531d2c8f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9bdac172";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7243337e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8ec9d585";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"613e3d82";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8bb6c783";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f3b1f75";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83cbcf90";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"7f3e2570";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65bfeba6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9a361d50";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58c6c7a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7403b3b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"30b1b4d3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6665645";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f8d9aba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb795035";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c8699bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd706a3a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a798ac6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d886772d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e6972b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"db9fa139";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1e4859bf";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c9b2b74d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3f2934a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bbd5d560";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5a2f2f83";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8fbecb81";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"70212c68";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88c4bf8c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8c3f375d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71c3d88c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d372f5f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5cabc4b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af46323e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4dbac1b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf514a31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b99b1cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc5f5b31";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3a8e98ca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ce7f6c33";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"388998c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d78b793b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e757dd1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd928739";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"285d73b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dcae9543";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"296e70cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e0a8b137";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"34494ab9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d2c3d251";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"403624a1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"afd9db7b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6835398f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9fcbdc7b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"7b3d3684";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92c5d177";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71422585";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83bbe080";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81402889";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88cde47c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a352673";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"64cce1a2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6371c68";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45c4d1ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5554254";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4dbbbaa7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b54b4e5e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3bb4b9ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b04f3e5e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41c6b1a7";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c8485153";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ab7b1b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b940533a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"30c394cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3596c34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"23a584d9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca678732";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e8575c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7728030";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41816ecc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b686943a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d7368cf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc899b22";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41644ecb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8a9ac32";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"43412ebf";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"9dc1cb5b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"67362da1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86cdc662";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"862d2a86";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6ec6c57b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8c333775";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"60d1bf96";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b373868";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"49d5b79d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ac2f4153";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40bab3ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ac354548";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44c4adb7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c9445f34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2caf95d5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c84a7327";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"2a9976cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd687d2d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"409183ca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb78882b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"377884cf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b77c822a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"49867ade";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d27c8b21";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"316b7dd2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3a7ad16";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"413e4cd4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0bcad2d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"53363db4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7cad14a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5d28509a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9ac4b465";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"692a3c93";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96c6b961";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68284495";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"91d8cb6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"722a3380";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9fd2d07c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74192d6a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"84d7db8d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74253861";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"73cfc29f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97343860";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75b8c89c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d403b56";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74becf97";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"963c3168";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74bbd89d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"99463655";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5dbceb9f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b93c2d53";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4eadc0b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5463d4b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42b1b7a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b45a4f50";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3facadb1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc414e4e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3da9a9ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d759633e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"27a89dc2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"da5d7938";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"33867ccc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d9739133";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f706eb6";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"d98cbc31";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"275b49b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0a1b952";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4f4a39a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aab8cd5e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5f4b3e99";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1add968";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6d45379a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2c0ca67";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74412a99";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74d5e982";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92362a89";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6cd3e491";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b931266c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4bc1cfa8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc483b4b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3fb8b3b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c25a5457";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48aca9ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3516150";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"46bbadaf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b84e4d49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"39b2a1cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d44f7233";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2bb196da";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e569952a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e906bd3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e1899b36";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"25695ec7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c296aa35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3f7659ca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b794a639";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"525b5ad1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"baa0a327";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b5f55d0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b6b9b538";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"524c41db";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b2c4c642";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"652e3eae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9fdad251";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5f333aac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96caba6e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6c3740a2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9cdbc05e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"71344098";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"99d8d072";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"66233396";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94e5c47f";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"77353479";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88f5ce98";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"89344476";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76c8c9a8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88322e62";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"69c1b3a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"89523a5d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65b5c3a6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"87403462";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fb0cc91";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b342853";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5cc4c9a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ad443840";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ea6c6cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb614739";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a9ea1c3";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"cd75662d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f7b98c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3797c4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c737fb2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d59b843e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"397f84ba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5909447";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"326567d2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"deacaf44";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"395a44a8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d4bfd953";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d3438aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adc9cb74";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"62352388";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9cdde07f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74403b7d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"84bed08c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"743e328c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8cbbcf85";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f412686";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81d7e587";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8f322b7f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61cbd495";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ac391e65";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50dad0a8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0504454";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3cacc3b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c9475a4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42b1a3b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca4c4253";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2dc6b5b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc4f5d47";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"2dae95c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d95b723e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2aad83c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd718840";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"219887cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d1718738";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"347f74d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d6878935";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3f7e78d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba899c3f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"428a77d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c27e7629";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"377b71d6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c9968825";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c6a72ee";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6aa9c34";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"475c59d8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bbac9a37";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"475754b1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2b3a657";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"435864b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfab8a50";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"465d6abf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2a8983d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"225c58c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"beb5ac4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b3b39af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c8bdbc54";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4440479c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1cdc16f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"563e3596";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9fbbbb79";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"664a3983";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"93b3cd64";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"584b3195";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"90b7cb7c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7e3a2182";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74cbde8c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"963e1f61";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"51bac99f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b046274a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38a5b3ce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c46b4f42";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"359faebc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb696240";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"378792bb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c3626351";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"349b9bbb";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"cb6c683b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"289183c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d47b8035";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"197463c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc84953f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"28775fbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c79aa043";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"356c5cb5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb87a43b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"416c4cc1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b498a331";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"406c49c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b49cc836";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"454a38c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7aac03a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50412fb4";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"92cecc49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"722d2ea1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"86c2d973";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8f2d2786";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"79bdbf6f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"81414582";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77c8bf78";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7932468d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8cbfc36f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7d202d79";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83e3cd7f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f1a3a72";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5fd9c3a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9e16364c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"60ccb699";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6314948";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"5ec4bbad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"90344554";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76bdc694";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8d433454";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7bbfd7a4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"95313d58";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5cbed3b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3423139";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58adc2a8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd4f423e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4299bfb9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3575547";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"52aba9ad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb5c4848";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3fa0baad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf52585a";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"33a6a4b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d95f5331";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"37989fc6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e36c7c30";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"247676cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d9869e3a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"376a60af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d7a1a548";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"356869b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c296b54e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"435747a8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4a9c448";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"57513a9f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a9b8db62";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5838369e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9cbfd470";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"743d1682";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7fd2da79";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8f343885";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6ebedc8f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a03a2c78";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6dbeba84";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"954b4875";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"67c7cf88";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"932c4481";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fd2c691";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ad322a6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"56e8d5a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc344a50";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45cab9c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca3c533f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45ba97bd";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"c2656f44";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31b89dc9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be596549";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ba393c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd58562e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"43b19ad5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba6a7727";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"349b93ec";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"da6c8220";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d7f7fd9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca8e8d1e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"396d7cdc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4969339";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50687acd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca987730";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b718dc0";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"ca8b8f38";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c6d7ecf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e79f8938";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"375b72ca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d9b1a330";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"285261bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cea4a452";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d5450b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ccaea654";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"456e6bae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b49f9e50";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c6747cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7a9a546";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"436342bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bdaec64b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e5641bb";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"a7afb85e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"545033b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a3c5c75f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"695543a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88b8c15b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"693e2ea5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8fb4ba6a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7443328c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ddacc6b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7c253281";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61c7c785";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a0192c64";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4bcabf96";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b441484e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2daea6b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc435545";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3aa18aac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b55d6a3f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"47a0a0ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7556d44";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"499d8fc6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca4d6624";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40a394d6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c869871d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38877ce4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d277931b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d716bd3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c494a02b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"426f67cc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b9a4a03e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"565f77d0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be9a9131";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"3d6a6fcc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c4a89c33";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d4663d7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cfc2b143";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a3256b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4d6ba46";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"553839aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a3d0bf6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"563d46a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2bec269";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"663e448c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4c5ba69";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"484347a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4c7d571";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5a3f2a97";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7d9dd78";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"6f3c2a7a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8fc0d283";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6d443989";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8ab9c975";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8344308c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83c1d37b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"833e2e92";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"75c7d685";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85492090";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7cd4c57b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88322e76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5dcece87";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9331397d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"58d1bd98";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b248386e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"56c3af9b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"873d5366";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5bbda39c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"973e3f60";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6cc8ba9c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97384455";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48ccb7b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b23b5136";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3fa89cd0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c65b6921";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3f9b8cd9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ba768c2a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e8169ca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b97b8c30";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"527274c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b38a9332";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"457083c9";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b98c8f25";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3f5a5dd3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c9a79c2f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41354fb8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"acc8c93e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"591c45a0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a4cec058";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"781f3f95";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97cabd71";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"74344387";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82d3b980";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6d323f85";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9ebcc578";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6d283672";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83ded582";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82302d63";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"76d7d7aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9d1b3043";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5dbfbfad";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a7464a33";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4db8b6b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a147444c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5baab8b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b34d3b36";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42adccb2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb58492f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"39a0aecd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb5c5741";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"328f98c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d4736628";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"218593c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d5776d3d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"296e83c8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d4848137";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"387782b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c97e7f3d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"218575c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d1667f38";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"228277c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e086981e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c7f60c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d18fa336";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"265642d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb8fa92d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e6d4eb2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b59dad3e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50586fbf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bf91a038";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"4a6b5fca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bca5aa20";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e4e58d4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfb8c63e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"602f47b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a1cccb41";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"682c3d9b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8cd8c16b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"85254695";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ccdbb70";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8f2d4473";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"84cac87f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"88333e7e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"76cec896";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9a21484d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6ad5c6a6";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"bb2c5538";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4bbdacbe";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c43e5e3b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3cab93da";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb666f26";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a968cc3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc6c8528";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"458285d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb757d43";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e8d89d3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb8c7f1b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"386689db";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c49b9e2b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e4e61db";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d0bca247";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"485959b9";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b9c9b548";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b3751b4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5b8ad58";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5b3f509f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bad0bb57";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54364da0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b6c9c369";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4436309e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfd0cc6a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"65322d88";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"94d5d885";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7720336c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"79d1d098";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"973e2b68";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"78c4d098";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8e4c4264";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"73b9d595";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8c3c2571";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"73c5c79b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"993b3176";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"56cbe194";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a63c215c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4bc1c7b0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c04a2b42";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ab2b4b0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc50534c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"35a9a8a3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af504d5f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ab0a7a9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c04a5750";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4bb7b7ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b53a5631";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"31b495c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d047693c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2fa587cf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d26e842a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d8c79c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb70862e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"46836acb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0818f36";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"458179be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be83972d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"397064d8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c58e8f28";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"465264ce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5aeb01c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"474251c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"acb3b252";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"5d3447af";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a9c5be4e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6541509d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"98c7ba64";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"69293da2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"97d0c373";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"80304081";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"83e3c97d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8228346c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"70dbc0a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a0274a62";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"67decdbb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b6395a2d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"46c6a0c9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc516836";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"479799d7";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b767633b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ea898c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b26c6a3f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3f97a0d8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0636234";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c8a8fde";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c791731c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d797fe5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc978529";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f606ed7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c8ab9834";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"365e5fc1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bfac924b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2e5f73c0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6969443";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"376463be";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"cda1913a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1f6047c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ccafbd4a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2a4646b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ccbcc049";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"444736aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4c9bf65";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"495141a7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9eb0be66";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"504f2faa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a9a7ac49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c5732b2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a4b9cf49";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4f352cb8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96cbc248";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"713516a0";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"84ccd963";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6e35388d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6fbbc274";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"862e2790";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ed3bb6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"79393f84";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"66cccb76";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8b213079";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6cc8b590";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9d303d5e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5cddc2a6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9e1f5244";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"46b9a8ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0304146";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"56bbb1b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ab4d5b39";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"4ba2abba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af595a44";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4f9c94bc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b655572f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4698a3cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6676b0c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f8693de";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d3847a1d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c636be4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6a3a81a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"464b5dbb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a8aeb043";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"544152b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2aea34e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"544d5ba7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b7c8ae48";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"4d3d51ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"abb5b557";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54243ea5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b1dad864";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5f262e72";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"96d6d47f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f192d6d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"77c9c69f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8a2a405f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7bc1d086";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7d45256a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7ab8d091";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7f363278";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"78bede8c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"962f2153";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6cc7dd8d";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"ab39245c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"49bbd4b3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5423754";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4cb5b1a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b55a4548";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"48a5b1a6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6464c63";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4cb6b4a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c83f394c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ac2acaa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8485649";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"28b4b4c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0425540";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"44b58eb3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c33f663e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"34b8a7c1";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"b1535d46";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4da59bc1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be48522d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4fa5a4c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a658661f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38a6a2dd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb546219";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3f8080ce";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c8767113";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2b748acb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b88a873c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"496771c6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c38b7941";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"42787baf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8898232";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2c7386cc";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"d99a893b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"374564c4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dbb4ac40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"353b54b1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1c2bf4b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4d4240a5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b5b7ba69";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61354e8a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aebcc369";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5d5b489e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"abbdc674";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5f43389f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"adbed57a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"593e1977";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"90d8ec8e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8e3d306e";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"70c6dcab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a5392a5d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5ec0d59c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aa553a5a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54b1c1ae";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a64f4a6a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"62b4af9f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0513a65";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4bd0c3a2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be43445d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"30c0c5c1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d6464f40";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"38b7a2c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c358604a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3fbda5be";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c04e7047";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"45b29cbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d2515f44";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"45bea7cc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb546c39";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3db6aad4";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ac5a5e2e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4f9c8cde";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c7646736";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c999ed3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2727633";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"449193d0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bb75613e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"54869fc1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd746440";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3aabaeb9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca5a5942";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"34969ed0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d7745f41";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1f8592cd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cd947b35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"32857bb9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca717b4d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b837cb3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b974774a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"34a189bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cc627e3a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2f8674db";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c6708225";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"31825ace";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c198a43c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"346c49c7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be97b24b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"475b53b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"afa1a73f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4e6a5aba";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a79d9c41";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4c5f56d1";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"af9ea633";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4b5247bb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b3c1ab3a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"443941bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a2ceb660";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5e293ea3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8dcdbd64";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7a39388c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7fd1b774";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"703a518e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"91bebb7e";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"7536387e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"87c7b67f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"892b3b60";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"61dad3ac";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"92303b57";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"5dc3b6bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ab403f3b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"56bea7b8";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9b564c45";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4ab6b3bf";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"a6503c4f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50ababb9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b4593d3d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"41acb3b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b0534449";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3ab1c1da";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"d755463c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"319e9aca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ce81662a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"199496c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c07a7152";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"40879bbc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c5725e46";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b9a99ab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc596146";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"20a993cc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"cb596f47";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2aa482ca";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e76e7b1d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"278e75dc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c084963d";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"337f66d8";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"be7e7e48";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"538e74bd";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bd797f35";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3c8e87cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b8716c2f";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"357f71ee";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca947d19";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"396c7bd2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"be9e9f30";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"375161cb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"b6a79445";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4d5862b9";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c0b8944b";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"396166b6";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"aab1964c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3d4551be";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"cabead52";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3e5447aa";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bbd8cf62";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"4a343e94";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9acec67a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"782d217e";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"8dd7ca88";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"6e404473";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"82bed493";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7e402f7a";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"7fc2beab";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"923b3863";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"68c6dea2";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"9d4a3853";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"50b7cdbe";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c2483c41";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------

Istart <= '1';
Iend <= '0';

Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Istart <= '0';
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"00000000";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"000088b5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;

Idata <= x"46a3a9c5";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"bc715c34";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3596a7cc";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"ca837641";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a7a86c3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d5867651";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3a7c83b0";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c998793c";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"2d7a8cc7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"dd898841";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"3b6e6ccb";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"e292ac32";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"1f664ec3";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"d9b9b849";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"384a40b7";
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
Idata <= x"c1baca5b";
Iend <= '1';
clk <= '1'; wait for 5 ns;
clk <= '0'; wait for 5 ns;
---------------------------------



Iend <= '0';

		
		  
		Ivalid <= '0';
		
		loop
		  clk <= '1'; wait for 5 ns;
		  clk <= '0'; wait for 5 ns;
        end loop;
      end process stimulus;
end architecture testbench; 
