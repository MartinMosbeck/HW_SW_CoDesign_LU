----------------------------------------------------------------------------------
-- Company:      TU Wien - ECS Group                                            --
-- Engineer:     Thomas Polzer                                                  --
--                                                                              --
-- Create Date:  21.09.2010                                                     --
-- Design Name:  DIDELU                                                         --
-- Module Name:  font_pkg                                                       --
-- Project Name: DIDELU                                                         --
-- Description:  Font ROM - Package - constant declaration of the font ROM.     --
--               The number of defined encodings, the character dimension       -- 
--               and the encoding itself are defiend in this package.           --
----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
--                                LIBRARIES                                     --
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.math_pkg.all;

----------------------------------------------------------------------------------
--                                 PACKAGE                                      --
----------------------------------------------------------------------------------

package font_pkg is
  constant CHAR_COUNT : integer := 256;
  constant CHAR_WIDTH : integer := 8;
  constant CHAR_HEIGHT : integer := 16;
 -- constant COLUMN_COUNT : integer := PIXEL_WIDTH / CHAR_WIDTH;
  --constant LINE_COUNT : integer := PIXEL_HEIGHT / CHAR_HEIGHT;
  type FONT_TYPE is array (0 to 2 ** (log2c(CHAR_COUNT) + log2c(CHAR_HEIGHT)) - 1) of std_logic_vector(0 to CHAR_WIDTH - 1);
 
 
	component font_rom is 
		port
		(
			vga_clk           : in std_logic;
			char              : in std_logic_vector(log2c(CHAR_COUNT) - 1 downto 0);
			char_height_pixel : in std_logic_vector(log2c(CHAR_HEIGHT) - 1 downto 0);
			decoded_char      : out std_logic_vector(0 to CHAR_WIDTH - 1)
		);
	end component;

 
 
  constant FONT_TABLE : FONT_TYPE :=
  (
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "10000001",
    "10100101",
    "10000001",
    "10000001",
    "10111101",
    "10011001",
    "10000001",
    "10000001",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "11111111",
    "11011011",
    "11111111",
    "11111111",
    "11000011",
    "11100111",
    "11111111",
    "11111111",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01101100",
    "11111110",
    "11111110",
    "11111110",
    "11111110",
    "01111100",
    "00111000",
    "00010000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00010000",
    "00111000",
    "01111100",
    "11111110",
    "01111100",
    "00111000",
    "00010000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00111100",
    "00111100",
    "11100111",
    "11100111",
    "11100111",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00111100",
    "01111110",
    "11111111",
    "11111111",
    "01111110",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00111100",
    "00111100",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11100111",
    "11000011",
    "11000011",
    "11100111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "01100110",
    "01000010",
    "01000010",
    "01100110",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11000011",
    "10011001",
    "10111101",
    "10111101",
    "10011001",
    "11000011",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00011110",
    "00001110",
    "00011010",
    "00110010",
    "01111000",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "01111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00111100",
    "00011000",
    "01111110",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111111",
    "00110011",
    "00111111",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "01110000",
    "11110000",
    "11100000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111111",
    "01100011",
    "01111111",
    "01100011",
    "01100011",
    "01100011",
    "01100011",
    "01100111",
    "11100111",
    "11100110",
    "11000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "11011011",
    "00111100",
    "11100111",
    "00111100",
    "11011011",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "10000000",
    "11000000",
    "11100000",
    "11110000",
    "11111000",
    "11111110",
    "11111000",
    "11110000",
    "11100000",
    "11000000",
    "10000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000010",
    "00000110",
    "00001110",
    "00011110",
    "00111110",
    "11111110",
    "00111110",
    "00011110",
    "00001110",
    "00000110",
    "00000010",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00111100",
    "01111110",
    "00011000",
    "00011000",
    "00011000",
    "01111110",
    "00111100",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00000000",
    "01100110",
    "01100110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111111",
    "11011011",
    "11011011",
    "11011011",
    "01111011",
    "00011011",
    "00011011",
    "00011011",
    "00011011",
    "00011011",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "01100000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "01101100",
    "00111000",
    "00001100",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "11111110",
    "11111110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00111100",
    "01111110",
    "00011000",
    "00011000",
    "00011000",
    "01111110",
    "00111100",
    "00011000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00111100",
    "01111110",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "01111110",
    "00111100",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00001100",
    "11111110",
    "00001100",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "01100000",
    "11111110",
    "01100000",
    "00110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000000",
    "11000000",
    "11000000",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00101000",
    "01101100",
    "11111110",
    "01101100",
    "00101000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00010000",
    "00111000",
    "00111000",
    "01111100",
    "01111100",
    "11111110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "11111110",
    "01111100",
    "01111100",
    "00111000",
    "00111000",
    "00010000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00111100",
    "00111100",
    "00111100",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "00100100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01101100",
    "01101100",
    "11111110",
    "01101100",
    "01101100",
    "01101100",
    "11111110",
    "01101100",
    "01101100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "01111100",
    "11000110",
    "11000010",
    "11000000",
    "01111100",
    "00000110",
    "00000110",
    "10000110",
    "11000110",
    "01111100",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000010",
    "11000110",
    "00001100",
    "00011000",
    "00110000",
    "01100000",
    "11000110",
    "10000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01101100",
    "01101100",
    "00111000",
    "01110110",
    "11011100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "00110000",
    "00110000",
    "01100000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001100",
    "00011000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00011000",
    "00001100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "00011000",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00011000",
    "00110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100110",
    "00111100",
    "11111111",
    "00111100",
    "01100110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "01111110",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000010",
    "00000110",
    "00001100",
    "00011000",
    "00110000",
    "01100000",
    "11000000",
    "10000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000", -- 0
    "00000000",	-- 1 
    "00000000",	-- 2
    "00111000",	-- 3
    "01101100",	-- 4
    "11000110", -- 5
    "11000110", -- 6
    "11010110", -- 7
    "11010110", -- 8
    "11000110", -- 9
    "11000110", -- A
    "01101100", -- B
    "00111000", -- C
    "00000000", -- D
    "00000000", -- E
    "00000000",	-- F
    "00000000", -- 0
    "00000000",	-- 1
    "00000000",	-- 2
    "00011000",	-- 3
    "00111000",	-- 4
    "01111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "00000110",
    "00001100",
    "00011000",
    "00110000",
    "01100000",
    "11000000",
    "11000110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "00000110",
    "00000110",
    "00111100",
    "00000110",
    "00000110",
    "00000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001100",
    "00011100",
    "00111100",
    "01101100",
    "11001100",
    "11111110",
    "00001100",
    "00001100",
    "00001100",
    "00011110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "11000000",
    "11000000",
    "11000000",
    "11111100",
    "00000110",
    "00000110",
    "00000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01100000",
    "11000000",
    "11000000",
    "11111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "11000110",
    "00000110",
    "00000110",
    "00001100",
    "00011000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "01111110",
    "00000110",
    "00000110",
    "00000110",
    "00001100",
    "01111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000110",
    "00001100",
    "00011000",
    "00110000",
    "01100000",
    "00110000",
    "00011000",
    "00001100",
    "00000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100000",
    "00110000",
    "00011000",
    "00001100",
    "00000110",
    "00001100",
    "00011000",
    "00110000",
    "01100000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "00001100",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11011110",
    "11011110",
    "11011110",
    "11011100",
    "11000000",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00010000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "11111110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111100",
    "01100110",
    "01100110",
    "01100110",
    "01111100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "11111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "01100110",
    "11000010",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000010",
    "01100110",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111000",
    "01101100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01101100",
    "11111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "01100110",
    "01100010",
    "01101000",
    "01111000",
    "01101000",
    "01100000",
    "01100010",
    "01100110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "01100110",
    "01100010",
    "01101000",
    "01111000",
    "01101000",
    "01100000",
    "01100000",
    "01100000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "01100110",
    "11000010",
    "11000000",
    "11000000",
    "11011110",
    "11000110",
    "11000110",
    "01100110",
    "00111010",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11111110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011110",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "11001100",
    "11001100",
    "11001100",
    "01111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11100110",
    "01100110",
    "01100110",
    "01101100",
    "01111000",
    "01111000",
    "01101100",
    "01100110",
    "01100110",
    "11100110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11110000",
    "01100000",
    "01100000",
    "01100000",
    "01100000",
    "01100000",
    "01100000",
    "01100010",
    "01100110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11101110",
    "11111110",
    "11111110",
    "11010110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11100110",
    "11110110",
    "11111110",
    "11011110",
    "11001110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111100",
    "01100110",
    "01100110",
    "01100110",
    "01111100",
    "01100000",
    "01100000",
    "01100000",
    "01100000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11010110",
    "11011110",
    "01111100",
    "00001100",
    "00001110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111100",
    "01100110",
    "01100110",
    "01100110",
    "01111100",
    "01101100",
    "01100110",
    "01100110",
    "01100110",
    "11100110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "01100000",
    "00111000",
    "00001100",
    "00000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "01111110",
    "01011010",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01101100",
    "00111000",
    "00010000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11010110",
    "11010110",
    "11010110",
    "11111110",
    "11101110",
    "01101100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11000110",
    "01101100",
    "01111100",
    "00111000",
    "00111000",
    "01111100",
    "01101100",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00111100",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "11000110",
    "10000110",
    "00001100",
    "00011000",
    "00110000",
    "01100000",
    "11000010",
    "11000110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "10000000",
    "11000000",
    "11100000",
    "01110000",
    "00111000",
    "00011100",
    "00001110",
    "00000110",
    "00000010",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00001100",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00010000",
    "00111000",
    "01101100",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "00011000",
    "00001100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111000",
    "00001100",
    "01111100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11100000",
    "01100000",
    "01100000",
    "01111000",
    "01101100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000000",
    "11000000",
    "11000000",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011100",
    "00001100",
    "00001100",
    "00111100",
    "01101100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11111110",
    "11000000",
    "11000000",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011100",
    "00110110",
    "00110010",
    "00110000",
    "01111000",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "01111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01110110",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "01111100",
    "00001100",
    "11001100",
    "01111000",
    "00000000",
    "00000000",
    "00000000",
    "11100000",
    "01100000",
    "01100000",
    "01101100",
    "01110110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "11100110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000110",
    "00000110",
    "00000000",
    "00001110",
    "00000110",
    "00000110",
    "00000110",
    "00000110",
    "00000110",
    "00000110",
    "01100110",
    "01100110",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "11100000",
    "01100000",
    "01100000",
    "01100110",
    "01101100",
    "01111000",
    "01111000",
    "01101100",
    "01100110",
    "11100110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11101100",
    "11111110",
    "11010110",
    "11010110",
    "11010110",
    "11010110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11011100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11011100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01111100",
    "01100000",
    "01100000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01110110",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "01111100",
    "00001100",
    "00001100",
    "00011110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11011100",
    "01110110",
    "01100110",
    "01100000",
    "01100000",
    "01100000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "01100000",
    "00111000",
    "00001100",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00010000",
    "00110000",
    "00110000",
    "11111100",
    "00110000",
    "00110000",
    "00110000",
    "00110000",
    "00110110",
    "00011100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01101100",
    "00111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11000110",
    "11010110",
    "11010110",
    "11010110",
    "11111110",
    "01101100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "01101100",
    "00111000",
    "00111000",
    "00111000",
    "01101100",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111110",
    "00000110",
    "00001100",
    "11111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "11001100",
    "00011000",
    "00110000",
    "01100000",
    "11000110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001110",
    "00011000",
    "00011000",
    "00011000",
    "01110000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00001110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01110000",
    "00011000",
    "00011000",
    "00011000",
    "00001110",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "01110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01110110",
    "11011100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00010000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "11000110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "01100110",
    "11000010",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000010",
    "01100110",
    "00111100",
    "00011000",
    "01110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11001100",
    "00000000",
    "00000000",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001100",
    "00011000",
    "00110000",
    "00000000",
    "01111100",
    "11000110",
    "11111110",
    "11000000",
    "11000000",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00010000",
    "00111000",
    "01101100",
    "00000000",
    "01111000",
    "00001100",
    "01111100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11001100",
    "00000000",
    "00000000",
    "01111000",
    "00001100",
    "01111100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100000",
    "00110000",
    "00011000",
    "00000000",
    "01111000",
    "00001100",
    "01111100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01101100",
    "00111000",
    "00000000",
    "01111000",
    "00001100",
    "01111100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000000",
    "11000000",
    "11000000",
    "11000110",
    "01111100",
    "00011000",
    "01110000",
    "00000000",
    "00000000",
    "00000000",
    "00010000",
    "00111000",
    "01101100",
    "00000000",
    "01111100",
    "11000110",
    "11111110",
    "11000000",
    "11000000",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11111110",
    "11000000",
    "11000000",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100000",
    "00110000",
    "00011000",
    "00000000",
    "01111100",
    "11000110",
    "11111110",
    "11000000",
    "11000000",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100110",
    "00000000",
    "00000000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00111100",
    "01100110",
    "00000000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100000",
    "00110000",
    "00011000",
    "00000000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "00000000",
    "00010000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "11111110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01101100",
    "00111000",
    "00010000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "11111110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001100",
    "00011000",
    "00000000",
    "11111110",
    "01100110",
    "01100010",
    "01101000",
    "01111000",
    "01101000",
    "01100010",
    "01100110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11101100",
    "00110110",
    "00110110",
    "01111110",
    "11011000",
    "11011000",
    "01101110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111110",
    "01101100",
    "11001100",
    "11001100",
    "11111110",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00010000",
    "00111000",
    "01101100",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100000",
    "00110000",
    "00011000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "01111000",
    "11001100",
    "00000000",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100000",
    "00110000",
    "00011000",
    "00000000",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "00000000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111110",
    "00000110",
    "00001100",
    "01111000",
    "00000000",
    "00000000",
    "11000110",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11001110",
    "11011110",
    "11110110",
    "11100110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01101100",
    "01100100",
    "01100000",
    "11110000",
    "01100000",
    "01100000",
    "01100000",
    "01100000",
    "11100110",
    "11111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000100",
    "01111100",
    "11001110",
    "11001110",
    "11010110",
    "11010110",
    "11010110",
    "11010110",
    "11100110",
    "11100110",
    "01111100",
    "01000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "01101100",
    "00111000",
    "00111000",
    "01101100",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001110",
    "00011011",
    "00011000",
    "00011000",
    "00011000",
    "01111110",
    "00011000",
    "00011000",
    "00011000",
    "11011000",
    "01110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00110000",
    "01100000",
    "00000000",
    "01111000",
    "00001100",
    "01111100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001100",
    "00011000",
    "00110000",
    "00000000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00110000",
    "01100000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00110000",
    "01100000",
    "00000000",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01110110",
    "11011100",
    "00000000",
    "11011100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01110110",
    "11011100",
    "00000000",
    "11000110",
    "11100110",
    "11110110",
    "11111110",
    "11011110",
    "11001110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "01101100",
    "01101100",
    "00111110",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01101100",
    "01101100",
    "00111000",
    "00000000",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "00110000",
    "00000000",
    "00110000",
    "00110000",
    "01100000",
    "11000000",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "10000010",
    "10110010",
    "10101010",
    "10110010",
    "10101010",
    "10101010",
    "10000010",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "00000110",
    "00000110",
    "00000110",
    "00000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100000",
    "11100000",
    "01100010",
    "01100110",
    "01101100",
    "00011000",
    "00110000",
    "01100000",
    "11011100",
    "10000110",
    "00001100",
    "00011000",
    "00111110",
    "00000000",
    "00000000",
    "00000000",
    "01100000",
    "11100000",
    "01100010",
    "01100110",
    "01101100",
    "00011000",
    "00110000",
    "01100110",
    "11001110",
    "10011010",
    "00111111",
    "00000110",
    "00000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00111100",
    "00111100",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110110",
    "01101100",
    "11011000",
    "01101100",
    "00110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11011000",
    "01101100",
    "00110110",
    "01101100",
    "11011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00010001",
    "01000100",
    "00010001",
    "01000100",
    "00010001",
    "01000100",
    "00010001",
    "01000100",
    "00010001",
    "01000100",
    "00010001",
    "01000100",
    "00010001",
    "01000100",
    "00010001",
    "01000100",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "11011101",
    "01110111",
    "11011101",
    "01110111",
    "11011101",
    "01110111",
    "11011101",
    "01110111",
    "11011101",
    "01110111",
    "11011101",
    "01110111",
    "11011101",
    "01110111",
    "11011101",
    "01110111",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "11111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "01100000",
    "11000000",
    "00010000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "11111110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "00010000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "11111110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001100",
    "00000110",
    "00010000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "11111110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "10000010",
    "10011010",
    "10100010",
    "10100010",
    "10100010",
    "10011010",
    "10000010",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "11110110",
    "00000110",
    "11110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "00000110",
    "11110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "11110110",
    "00000110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "01111100",
    "11000110",
    "11000000",
    "11000000",
    "11000110",
    "01111100",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100110",
    "01100110",
    "00111100",
    "00011000",
    "01111110",
    "00011000",
    "01111110",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011111",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "11111111",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "01110110",
    "11011100",
    "00000000",
    "01111000",
    "00001100",
    "01111100",
    "11001100",
    "11001100",
    "11001100",
    "01110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01110110",
    "11011100",
    "00000000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "11111110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110111",
    "00110000",
    "00111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111111",
    "00110000",
    "00110111",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "11110111",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "11110111",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110111",
    "00110000",
    "00110111",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "11110111",
    "00000000",
    "11110111",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00110110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110100",
    "00011000",
    "00101100",
    "00000110",
    "00111110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111000",
    "01101100",
    "01100110",
    "01100110",
    "11110110",
    "01100110",
    "01100110",
    "01100110",
    "01101100",
    "11111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01101100",
    "00000000",
    "11111110",
    "01100110",
    "01100010",
    "01101000",
    "01111000",
    "01101000",
    "01100010",
    "01100110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "00000000",
    "11111110",
    "01100110",
    "01100010",
    "01101000",
    "01111000",
    "01101000",
    "01100010",
    "01100110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "00011000",
    "00000000",
    "11111110",
    "01100110",
    "01100010",
    "01101000",
    "01111000",
    "01101000",
    "01100010",
    "01100110",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001100",
    "00011000",
    "00000000",
    "00111100",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "01100110",
    "00000000",
    "00111100",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100110",
    "00000000",
    "00111100",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "11111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011111",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "00011000",
    "00000000",
    "00111100",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00110000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111000",
    "11001100",
    "11001100",
    "11001100",
    "11011000",
    "11001100",
    "11000110",
    "11000110",
    "11000110",
    "11001100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01101100",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "00011000",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01110110",
    "11011100",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01110110",
    "11011100",
    "00000000",
    "01111100",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01111100",
    "01100000",
    "01100000",
    "11000000",
    "00000000",
    "00000000",
    "00000000",
    "11100000",
    "01100000",
    "01100000",
    "01111100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01111100",
    "01100000",
    "01100000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "11110000",
    "01100000",
    "01111100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01111100",
    "01100000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00110000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01101100",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00110000",
    "00011000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001100",
    "00011000",
    "00110000",
    "00000000",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "11000110",
    "01111110",
    "00000110",
    "00001100",
    "11111000",
    "00000000",
    "00001100",
    "00011000",
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00111100",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001100",
    "00011000",
    "00110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "01111110",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "11100000",
    "00110000",
    "01100010",
    "00110110",
    "11101100",
    "00011000",
    "00110000",
    "01100110",
    "11001110",
    "10011010",
    "00111111",
    "00000110",
    "00000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111111",
    "11011011",
    "11011011",
    "11011011",
    "01111011",
    "00011011",
    "00011011",
    "00011011",
    "00011011",
    "00011011",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "11000110",
    "01100000",
    "00111000",
    "01101100",
    "11000110",
    "11000110",
    "01101100",
    "00111000",
    "00001100",
    "11000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00000000",
    "01111110",
    "00000000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00001100",
    "01111000",
    "00000000",
    "00000000",
    "00000000",
    "00111000",
    "01101100",
    "01101100",
    "00111000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11000110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111100",
    "00000110",
    "00111100",
    "00000110",
    "00000110",
    "01111100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111100",
    "01100110",
    "00001100",
    "00011000",
    "00110010",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "01111110",
    "01111110",
    "01111110",
    "01111110",
    "01111110",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000"
  );
end package font_pkg;

--- EOF ---
