library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.audiocore_pkg.all;

entity outputlogic is
	port 
	(
		clk : in std_logic;
		res_n : in std_logic;

		data_in : in fixpoint;
		validin : in std_logic;
		
		data_out : out byte;
		validout : out std_logic
	);
end outputlogic;

architecture behavior of outputlogic is
	signal data_out_cur,data_out_next : byte; 
	signal data : fixpoint;
	signal validout_cur, validout_next, valid : std_logic;

	function fixpoint_mult(a,b:fixpoint) return fixpoint is
				variable result_full : fixpoint_product;
	begin
		result_full := a * b;

		return result_full(55 downto 24);
	end function;
begin

	deci: decimator
	generic map
	(
		N => 2
	)	
	port map 
	(
		clk =>clk,
		res_n =>res_n,

		data_in =>data_in,
		validin =>validin,
		
		data_out =>data, 
		validout => valid
	);


	do_output: process (data,valid)
		constant factor : fixpoint := x"1e000000";
		variable data_fixp : fixpoint;
		constant v127 : signed(7 downto 0) := "01111111"; 
		
		variable factor0 : fixpoint;
		variable product : fixpoint_product;
	begin
		data_out_next <= data_out_cur;
		validout_next <= validout_cur;

		if(valid = '0') then
			validout_next <= '0';
		else
			validout_next <= '1';
			
			--sign extend
--			if(data(31) = '1' then
--				factor0(63 downto 56) := (others => '1');
--			else
--				factor0(63 downto 56) := (others => '0');
--			end if;
--			factor0(23 downto 0) := (others => '0');
--			factor0(55 downto 24) := data;
--
--			factor1(63 downto 48) := to_signed(30, 16);
--			factor1(47 downto 0) := (others => '0');
--			product := factor0 * factor1;
--			data_out_next <= product(103 downto 71);

			data_fixp := fixpoint_mult(data,factor);
			data_out_next <= std_logic_vector(data_fixp(31 downto 24) + v127);
			
		end if; 
	end process do_output;

	sync: process (clk,res_n)
	begin
		if res_n = '0' then
			data_out_cur <= (others =>'0');
			validout_cur <= '0';
		elsif rising_edge(clk) then
			--internals
				data_out_cur <= data_out_next;
				validout_cur <= validout_next;
			--outputs
				data_out <= data_out_next;
				validout <= validout_next;
		end if;
	end process sync;

end behavior;
