
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package audiocore_pkg is
	subtype fixedpoint is signed(31 downto 0);
	subtype byte is std_logic_vector(7 downto 0);
	subtype sgdma_frame is std_logic_vector(31 downto 0);
	subtype index_time is integer range 0 to 24; 
end package audiocore_pkg;

package body audiocore_pkg is

	function lookup_sin(index:index_time) 
		return fixedpoint is
	begin 
		case index is
			when 0 =>
				return "10000000000000000000000000000000";
			when 1 =>
				return "00000000111111110111111010101101";
			when 2 =>
				return "00000000001000000001010111010110";
			when 3 =>
				return "10000000111110110111011100101101";
			when 4 =>
				return "10000000001111111010101000100011";
			when 5 =>
				return "00000000111100110111100001110000";
			when 6 =>
				return "00000000010111100011110101101001";
			when 7 =>
				return "10000000111001111010001010111110";
			when 8 =>
				return "10000000011110110101010000110101";
			when 9 =>
				return "00000000110110000010010111011111";
			when 10 =>
				return "00000000100101100111100100011000";
			when 11 =>
				return "10000000110001010100000001011011";
			when 12 =>
				return "10000000101011110011111001111010";
			when 13 =>
				return "00000000101011110011111001111010";
			when 14 =>
				return "00000000110001010100000001011011";
			when 15 =>
				return "10000000100101100111100100011000";
			when 16 =>
				return "10000000110110000010010111011111";
			when 17 =>
				return "00000000011110110101010000110101";
			when 18 =>
				return "00000000111001111010001010111110";
			when 19 =>
				return "10000000010111100011110101101001";
			when 20 =>
				return "10000000111100110111100001110000";
			when 21 =>
				return "00000000001111111010101000100011";
			when 22 =>
				return "00000000111110110111011100101101";
			when 23 =>
				return "10000000001000000001010111010110";
			when 24 =>
				return "10000000111111110111111010101101";
		end case;
	end function;

	function lookup_cos(index:index_time)
		return fixedpoint is
	begin	
		case index is
			when 0 =>
				return "00000001000000000000000000000000";
			when 1 =>
				return "00000000000100000001001100001010";
			when 2 =>
				return "10000000111111011111101100111010";
			when 3 =>
				return "10000000001011111111100000111000";
			when 4 =>
				return "00000000111101111111010100010000";
			when 5 =>
				return "00000000010011110001101110111100";
			when 6 =>
				return "10000000111011100000010111010100";
			when 7 =>
				return "10000000011011001111111111011111";
			when 8 =>
				return "00000000111000000101010110100010";
			when 9 =>
				return "00000000100010010010101111110001";
			when 10 =>
				return "10000000110011110001101110111100";
			when 11 =>
				return "10000000101000110010111000110111";
			when 12 =>
				return "00000000101110101001110110110000";
			when 13 =>
				return "00000000101110101001110110110000";
			when 14 =>
				return "10000000101000110010111000110111";
			when 15 =>
				return "10000000110011110001101110111100";
			when 16 =>
				return "00000000100010010010101111110001";
			when 17 =>
				return "00000000111000000101010110100010";
			when 18 =>
				return "10000000011011001111111111011111";
			when 19 =>
				return "10000000111011100000010111010100";
			when 20 =>
				return "00000000010011110001101110111100";
			when 21 =>
				return "00000000111101111111010100010000";
			when 22 =>
				return "10000000001011111111100000111000";
			when 23 =>
				return "10000000111111011111101100111010";
			when 24 =>
				return "00000000000100000001001100001010";
		end case;
	end function;

end package body;


